
`include "dump_file_agent.svh"
`include "csv_file_dump.svh"
`include "sample_agent.svh"
`include "loop_sample_agent.svh"
`include "sample_manager.svh"
`include "nodf_module_interface.svh"
`include "nodf_module_monitor.svh"
`include "seq_loop_interface.svh"
`include "seq_loop_monitor.svh"
`include "upc_loop_interface.svh"
`include "upc_loop_monitor.svh"
`timescale 1ns/1ps

// top module for dataflow related monitors
module dataflow_monitor(
input logic clock,
input logic reset,
input logic finish
);



    nodf_module_intf module_intf_1(clock,reset);
    assign module_intf_1.ap_start = AESL_inst_master.ap_start;
    assign module_intf_1.ap_ready = AESL_inst_master.ap_ready;
    assign module_intf_1.ap_done = AESL_inst_master.ap_done;
    assign module_intf_1.ap_continue = 1'b1;
    assign module_intf_1.finish = finish;
    csv_file_dump mstatus_csv_dumper_1;
    nodf_module_monitor module_monitor_1;
    nodf_module_intf module_intf_2(clock,reset);
    assign module_intf_2.ap_start = AESL_inst_master.grp_convolution1_1_fu_326.ap_start;
    assign module_intf_2.ap_ready = AESL_inst_master.grp_convolution1_1_fu_326.ap_ready;
    assign module_intf_2.ap_done = AESL_inst_master.grp_convolution1_1_fu_326.ap_done;
    assign module_intf_2.ap_continue = 1'b1;
    assign module_intf_2.finish = finish;
    csv_file_dump mstatus_csv_dumper_2;
    nodf_module_monitor module_monitor_2;
    nodf_module_intf module_intf_3(clock,reset);
    assign module_intf_3.ap_start = AESL_inst_master.grp_maxPool_1_fu_338.ap_start;
    assign module_intf_3.ap_ready = AESL_inst_master.grp_maxPool_1_fu_338.ap_ready;
    assign module_intf_3.ap_done = AESL_inst_master.grp_maxPool_1_fu_338.ap_done;
    assign module_intf_3.ap_continue = 1'b1;
    assign module_intf_3.finish = finish;
    csv_file_dump mstatus_csv_dumper_3;
    nodf_module_monitor module_monitor_3;
    nodf_module_intf module_intf_4(clock,reset);
    assign module_intf_4.ap_start = AESL_inst_master.grp_convolution2_fu_344.ap_start;
    assign module_intf_4.ap_ready = AESL_inst_master.grp_convolution2_fu_344.ap_ready;
    assign module_intf_4.ap_done = AESL_inst_master.grp_convolution2_fu_344.ap_done;
    assign module_intf_4.ap_continue = 1'b1;
    assign module_intf_4.finish = finish;
    csv_file_dump mstatus_csv_dumper_4;
    nodf_module_monitor module_monitor_4;
    nodf_module_intf module_intf_5(clock,reset);
    assign module_intf_5.ap_start = AESL_inst_master.grp_maxPool_fu_354.ap_start;
    assign module_intf_5.ap_ready = AESL_inst_master.grp_maxPool_fu_354.ap_ready;
    assign module_intf_5.ap_done = AESL_inst_master.grp_maxPool_fu_354.ap_done;
    assign module_intf_5.ap_continue = 1'b1;
    assign module_intf_5.finish = finish;
    csv_file_dump mstatus_csv_dumper_5;
    nodf_module_monitor module_monitor_5;
    nodf_module_intf module_intf_6(clock,reset);
    assign module_intf_6.ap_start = AESL_inst_master.grp_master_Pipeline_VITIS_LOOP_143_2_fu_360.ap_start;
    assign module_intf_6.ap_ready = AESL_inst_master.grp_master_Pipeline_VITIS_LOOP_143_2_fu_360.ap_ready;
    assign module_intf_6.ap_done = AESL_inst_master.grp_master_Pipeline_VITIS_LOOP_143_2_fu_360.ap_done;
    assign module_intf_6.ap_continue = 1'b1;
    assign module_intf_6.finish = finish;
    csv_file_dump mstatus_csv_dumper_6;
    nodf_module_monitor module_monitor_6;

    seq_loop_intf#(48) seq_loop_intf_1(clock,reset);
    assign seq_loop_intf_1.pre_loop_state0 = AESL_inst_master.ap_ST_fsm_state11;
    assign seq_loop_intf_1.pre_states_valid = 1'b1;
    assign seq_loop_intf_1.post_loop_state0 = AESL_inst_master.ap_ST_fsm_state11;
    assign seq_loop_intf_1.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_1.post_loop_state1 = 48'h0;
    assign seq_loop_intf_1.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_1.post_loop_state2 = 48'h0;
    assign seq_loop_intf_1.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_1.quit_loop_state0 = AESL_inst_master.ap_ST_fsm_state12;
    assign seq_loop_intf_1.quit_states_valid = 1'b1;
    assign seq_loop_intf_1.cur_state = AESL_inst_master.ap_CS_fsm;
    assign seq_loop_intf_1.iter_start_state = AESL_inst_master.ap_ST_fsm_state12;
    assign seq_loop_intf_1.iter_end_state0 = AESL_inst_master.ap_ST_fsm_state19;
    assign seq_loop_intf_1.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_1.one_state_loop = 1'b0;
    assign seq_loop_intf_1.one_state_block = 1'b0;
    assign seq_loop_intf_1.finish = finish;
    csv_file_dump seq_loop_csv_dumper_1;
    seq_loop_monitor #(48) seq_loop_monitor_1;
    seq_loop_intf#(48) seq_loop_intf_2(clock,reset);
    assign seq_loop_intf_2.pre_loop_state0 = AESL_inst_master.ap_ST_fsm_state10;
    assign seq_loop_intf_2.pre_states_valid = 1'b1;
    assign seq_loop_intf_2.post_loop_state0 = AESL_inst_master.ap_ST_fsm_state20;
    assign seq_loop_intf_2.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_2.post_loop_state1 = 48'h0;
    assign seq_loop_intf_2.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_2.post_loop_state2 = 48'h0;
    assign seq_loop_intf_2.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_2.quit_loop_state0 = AESL_inst_master.ap_ST_fsm_state11;
    assign seq_loop_intf_2.quit_states_valid = 1'b1;
    assign seq_loop_intf_2.cur_state = AESL_inst_master.ap_CS_fsm;
    assign seq_loop_intf_2.iter_start_state = AESL_inst_master.ap_ST_fsm_state11;
    assign seq_loop_intf_2.iter_end_state0 = AESL_inst_master.ap_ST_fsm_state12;
    assign seq_loop_intf_2.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_2.one_state_loop = 1'b0;
    assign seq_loop_intf_2.one_state_block = 1'b0;
    assign seq_loop_intf_2.finish = finish;
    csv_file_dump seq_loop_csv_dumper_2;
    seq_loop_monitor #(48) seq_loop_monitor_2;
    seq_loop_intf#(48) seq_loop_intf_3(clock,reset);
    assign seq_loop_intf_3.pre_loop_state0 = AESL_inst_master.ap_ST_fsm_state8;
    assign seq_loop_intf_3.pre_states_valid = 1'b1;
    assign seq_loop_intf_3.post_loop_state0 = AESL_inst_master.ap_ST_fsm_state21;
    assign seq_loop_intf_3.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_3.post_loop_state1 = 48'h0;
    assign seq_loop_intf_3.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_3.post_loop_state2 = 48'h0;
    assign seq_loop_intf_3.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_3.quit_loop_state0 = AESL_inst_master.ap_ST_fsm_state9;
    assign seq_loop_intf_3.quit_states_valid = 1'b1;
    assign seq_loop_intf_3.cur_state = AESL_inst_master.ap_CS_fsm;
    assign seq_loop_intf_3.iter_start_state = AESL_inst_master.ap_ST_fsm_state9;
    assign seq_loop_intf_3.iter_end_state0 = AESL_inst_master.ap_ST_fsm_state20;
    assign seq_loop_intf_3.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_3.one_state_loop = 1'b0;
    assign seq_loop_intf_3.one_state_block = 1'b0;
    assign seq_loop_intf_3.finish = finish;
    csv_file_dump seq_loop_csv_dumper_3;
    seq_loop_monitor #(48) seq_loop_monitor_3;
    seq_loop_intf#(48) seq_loop_intf_4(clock,reset);
    assign seq_loop_intf_4.pre_loop_state0 = AESL_inst_master.ap_ST_fsm_state21;
    assign seq_loop_intf_4.pre_states_valid = 1'b1;
    assign seq_loop_intf_4.post_loop_state0 = AESL_inst_master.ap_ST_fsm_state21;
    assign seq_loop_intf_4.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_4.post_loop_state1 = 48'h0;
    assign seq_loop_intf_4.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_4.post_loop_state2 = 48'h0;
    assign seq_loop_intf_4.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_4.quit_loop_state0 = AESL_inst_master.ap_ST_fsm_state22;
    assign seq_loop_intf_4.quit_states_valid = 1'b1;
    assign seq_loop_intf_4.cur_state = AESL_inst_master.ap_CS_fsm;
    assign seq_loop_intf_4.iter_start_state = AESL_inst_master.ap_ST_fsm_state22;
    assign seq_loop_intf_4.iter_end_state0 = AESL_inst_master.ap_ST_fsm_state29;
    assign seq_loop_intf_4.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_4.one_state_loop = 1'b0;
    assign seq_loop_intf_4.one_state_block = 1'b0;
    assign seq_loop_intf_4.finish = finish;
    csv_file_dump seq_loop_csv_dumper_4;
    seq_loop_monitor #(48) seq_loop_monitor_4;
    seq_loop_intf#(48) seq_loop_intf_5(clock,reset);
    assign seq_loop_intf_5.pre_loop_state0 = AESL_inst_master.ap_ST_fsm_state9;
    assign seq_loop_intf_5.pre_states_valid = 1'b1;
    assign seq_loop_intf_5.post_loop_state0 = AESL_inst_master.ap_ST_fsm_state30;
    assign seq_loop_intf_5.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_5.post_loop_state1 = 48'h0;
    assign seq_loop_intf_5.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_5.post_loop_state2 = 48'h0;
    assign seq_loop_intf_5.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_5.quit_loop_state0 = AESL_inst_master.ap_ST_fsm_state21;
    assign seq_loop_intf_5.quit_states_valid = 1'b1;
    assign seq_loop_intf_5.cur_state = AESL_inst_master.ap_CS_fsm;
    assign seq_loop_intf_5.iter_start_state = AESL_inst_master.ap_ST_fsm_state21;
    assign seq_loop_intf_5.iter_end_state0 = AESL_inst_master.ap_ST_fsm_state22;
    assign seq_loop_intf_5.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_5.one_state_loop = 1'b0;
    assign seq_loop_intf_5.one_state_block = 1'b0;
    assign seq_loop_intf_5.finish = finish;
    csv_file_dump seq_loop_csv_dumper_5;
    seq_loop_monitor #(48) seq_loop_monitor_5;
    seq_loop_intf#(48) seq_loop_intf_6(clock,reset);
    assign seq_loop_intf_6.pre_loop_state0 = AESL_inst_master.ap_ST_fsm_state21;
    assign seq_loop_intf_6.pre_states_valid = 1'b1;
    assign seq_loop_intf_6.post_loop_state0 = AESL_inst_master.ap_ST_fsm_state48;
    assign seq_loop_intf_6.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_6.post_loop_state1 = 48'h0;
    assign seq_loop_intf_6.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_6.post_loop_state2 = 48'h0;
    assign seq_loop_intf_6.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_6.quit_loop_state0 = AESL_inst_master.ap_ST_fsm_state30;
    assign seq_loop_intf_6.quit_states_valid = 1'b1;
    assign seq_loop_intf_6.cur_state = AESL_inst_master.ap_CS_fsm;
    assign seq_loop_intf_6.iter_start_state = AESL_inst_master.ap_ST_fsm_state30;
    assign seq_loop_intf_6.iter_end_state0 = AESL_inst_master.ap_ST_fsm_state47;
    assign seq_loop_intf_6.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_6.one_state_loop = 1'b0;
    assign seq_loop_intf_6.one_state_block = 1'b0;
    assign seq_loop_intf_6.finish = finish;
    csv_file_dump seq_loop_csv_dumper_6;
    seq_loop_monitor #(48) seq_loop_monitor_6;
    seq_loop_intf#(130) seq_loop_intf_7(clock,reset);
    assign seq_loop_intf_7.pre_loop_state0 = AESL_inst_master.grp_convolution1_1_fu_326.ap_ST_fsm_state4;
    assign seq_loop_intf_7.pre_states_valid = 1'b1;
    assign seq_loop_intf_7.post_loop_state0 = AESL_inst_master.grp_convolution1_1_fu_326.ap_ST_fsm_state4;
    assign seq_loop_intf_7.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_7.post_loop_state1 = 130'h0;
    assign seq_loop_intf_7.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_7.post_loop_state2 = 130'h0;
    assign seq_loop_intf_7.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_7.quit_loop_state0 = AESL_inst_master.grp_convolution1_1_fu_326.ap_ST_fsm_state5;
    assign seq_loop_intf_7.quit_states_valid = 1'b1;
    assign seq_loop_intf_7.cur_state = AESL_inst_master.grp_convolution1_1_fu_326.ap_CS_fsm;
    assign seq_loop_intf_7.iter_start_state = AESL_inst_master.grp_convolution1_1_fu_326.ap_ST_fsm_state5;
    assign seq_loop_intf_7.iter_end_state0 = AESL_inst_master.grp_convolution1_1_fu_326.ap_ST_fsm_state130;
    assign seq_loop_intf_7.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_7.one_state_loop = 1'b0;
    assign seq_loop_intf_7.one_state_block = 1'b0;
    assign seq_loop_intf_7.finish = finish;
    csv_file_dump seq_loop_csv_dumper_7;
    seq_loop_monitor #(130) seq_loop_monitor_7;
    seq_loop_intf#(130) seq_loop_intf_8(clock,reset);
    assign seq_loop_intf_8.pre_loop_state0 = AESL_inst_master.grp_convolution1_1_fu_326.ap_ST_fsm_state3;
    assign seq_loop_intf_8.pre_states_valid = 1'b1;
    assign seq_loop_intf_8.post_loop_state0 = AESL_inst_master.grp_convolution1_1_fu_326.ap_ST_fsm_state2;
    assign seq_loop_intf_8.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_8.post_loop_state1 = 130'h0;
    assign seq_loop_intf_8.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_8.post_loop_state2 = 130'h0;
    assign seq_loop_intf_8.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_8.quit_loop_state0 = AESL_inst_master.grp_convolution1_1_fu_326.ap_ST_fsm_state4;
    assign seq_loop_intf_8.quit_states_valid = 1'b1;
    assign seq_loop_intf_8.cur_state = AESL_inst_master.grp_convolution1_1_fu_326.ap_CS_fsm;
    assign seq_loop_intf_8.iter_start_state = AESL_inst_master.grp_convolution1_1_fu_326.ap_ST_fsm_state4;
    assign seq_loop_intf_8.iter_end_state0 = AESL_inst_master.grp_convolution1_1_fu_326.ap_ST_fsm_state5;
    assign seq_loop_intf_8.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_8.one_state_loop = 1'b0;
    assign seq_loop_intf_8.one_state_block = 1'b0;
    assign seq_loop_intf_8.finish = finish;
    csv_file_dump seq_loop_csv_dumper_8;
    seq_loop_monitor #(130) seq_loop_monitor_8;
    seq_loop_intf#(130) seq_loop_intf_9(clock,reset);
    assign seq_loop_intf_9.pre_loop_state0 = AESL_inst_master.grp_convolution1_1_fu_326.ap_ST_fsm_state1;
    assign seq_loop_intf_9.pre_states_valid = 1'b1;
    assign seq_loop_intf_9.post_loop_state0 = AESL_inst_master.grp_convolution1_1_fu_326.ap_ST_fsm_state1;
    assign seq_loop_intf_9.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_9.post_loop_state1 = 130'h0;
    assign seq_loop_intf_9.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_9.post_loop_state2 = 130'h0;
    assign seq_loop_intf_9.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_9.quit_loop_state0 = AESL_inst_master.grp_convolution1_1_fu_326.ap_ST_fsm_state2;
    assign seq_loop_intf_9.quit_states_valid = 1'b1;
    assign seq_loop_intf_9.cur_state = AESL_inst_master.grp_convolution1_1_fu_326.ap_CS_fsm;
    assign seq_loop_intf_9.iter_start_state = AESL_inst_master.grp_convolution1_1_fu_326.ap_ST_fsm_state2;
    assign seq_loop_intf_9.iter_end_state0 = AESL_inst_master.grp_convolution1_1_fu_326.ap_ST_fsm_state4;
    assign seq_loop_intf_9.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_9.one_state_loop = 1'b0;
    assign seq_loop_intf_9.one_state_block = 1'b0;
    assign seq_loop_intf_9.finish = finish;
    csv_file_dump seq_loop_csv_dumper_9;
    seq_loop_monitor #(130) seq_loop_monitor_9;
    seq_loop_intf#(20) seq_loop_intf_10(clock,reset);
    assign seq_loop_intf_10.pre_loop_state0 = AESL_inst_master.grp_maxPool_1_fu_338.ap_ST_fsm_state15;
    assign seq_loop_intf_10.pre_states_valid = 1'b1;
    assign seq_loop_intf_10.post_loop_state0 = AESL_inst_master.grp_maxPool_1_fu_338.ap_ST_fsm_state3;
    assign seq_loop_intf_10.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_10.post_loop_state1 = 20'h0;
    assign seq_loop_intf_10.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_10.post_loop_state2 = 20'h0;
    assign seq_loop_intf_10.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_10.quit_loop_state0 = AESL_inst_master.grp_maxPool_1_fu_338.ap_ST_fsm_state16;
    assign seq_loop_intf_10.quit_states_valid = 1'b1;
    assign seq_loop_intf_10.cur_state = AESL_inst_master.grp_maxPool_1_fu_338.ap_CS_fsm;
    assign seq_loop_intf_10.iter_start_state = AESL_inst_master.grp_maxPool_1_fu_338.ap_ST_fsm_state16;
    assign seq_loop_intf_10.iter_end_state0 = AESL_inst_master.grp_maxPool_1_fu_338.ap_ST_fsm_state20;
    assign seq_loop_intf_10.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_10.one_state_loop = 1'b0;
    assign seq_loop_intf_10.one_state_block = 1'b0;
    assign seq_loop_intf_10.finish = finish;
    csv_file_dump seq_loop_csv_dumper_10;
    seq_loop_monitor #(20) seq_loop_monitor_10;
    seq_loop_intf#(20) seq_loop_intf_11(clock,reset);
    assign seq_loop_intf_11.pre_loop_state0 = AESL_inst_master.grp_maxPool_1_fu_338.ap_ST_fsm_state2;
    assign seq_loop_intf_11.pre_states_valid = 1'b1;
    assign seq_loop_intf_11.post_loop_state0 = AESL_inst_master.grp_maxPool_1_fu_338.ap_ST_fsm_state2;
    assign seq_loop_intf_11.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_11.post_loop_state1 = 20'h0;
    assign seq_loop_intf_11.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_11.post_loop_state2 = 20'h0;
    assign seq_loop_intf_11.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_11.quit_loop_state0 = AESL_inst_master.grp_maxPool_1_fu_338.ap_ST_fsm_state3;
    assign seq_loop_intf_11.quit_states_valid = 1'b1;
    assign seq_loop_intf_11.cur_state = AESL_inst_master.grp_maxPool_1_fu_338.ap_CS_fsm;
    assign seq_loop_intf_11.iter_start_state = AESL_inst_master.grp_maxPool_1_fu_338.ap_ST_fsm_state3;
    assign seq_loop_intf_11.iter_end_state0 = AESL_inst_master.grp_maxPool_1_fu_338.ap_ST_fsm_state16;
    assign seq_loop_intf_11.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_11.one_state_loop = 1'b0;
    assign seq_loop_intf_11.one_state_block = 1'b0;
    assign seq_loop_intf_11.finish = finish;
    csv_file_dump seq_loop_csv_dumper_11;
    seq_loop_monitor #(20) seq_loop_monitor_11;
    seq_loop_intf#(20) seq_loop_intf_12(clock,reset);
    assign seq_loop_intf_12.pre_loop_state0 = AESL_inst_master.grp_maxPool_1_fu_338.ap_ST_fsm_state1;
    assign seq_loop_intf_12.pre_states_valid = 1'b1;
    assign seq_loop_intf_12.post_loop_state0 = AESL_inst_master.grp_maxPool_1_fu_338.ap_ST_fsm_state1;
    assign seq_loop_intf_12.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_12.post_loop_state1 = 20'h0;
    assign seq_loop_intf_12.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_12.post_loop_state2 = 20'h0;
    assign seq_loop_intf_12.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_12.quit_loop_state0 = AESL_inst_master.grp_maxPool_1_fu_338.ap_ST_fsm_state2;
    assign seq_loop_intf_12.quit_states_valid = 1'b1;
    assign seq_loop_intf_12.cur_state = AESL_inst_master.grp_maxPool_1_fu_338.ap_CS_fsm;
    assign seq_loop_intf_12.iter_start_state = AESL_inst_master.grp_maxPool_1_fu_338.ap_ST_fsm_state2;
    assign seq_loop_intf_12.iter_end_state0 = AESL_inst_master.grp_maxPool_1_fu_338.ap_ST_fsm_state3;
    assign seq_loop_intf_12.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_12.one_state_loop = 1'b0;
    assign seq_loop_intf_12.one_state_block = 1'b0;
    assign seq_loop_intf_12.finish = finish;
    csv_file_dump seq_loop_csv_dumper_12;
    seq_loop_monitor #(20) seq_loop_monitor_12;
    seq_loop_intf#(42) seq_loop_intf_13(clock,reset);
    assign seq_loop_intf_13.pre_loop_state0 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state4;
    assign seq_loop_intf_13.pre_states_valid = 1'b1;
    assign seq_loop_intf_13.post_loop_state0 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state13;
    assign seq_loop_intf_13.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_13.post_loop_state1 = 42'h0;
    assign seq_loop_intf_13.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_13.post_loop_state2 = 42'h0;
    assign seq_loop_intf_13.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_13.quit_loop_state0 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state5;
    assign seq_loop_intf_13.quit_states_valid = 1'b1;
    assign seq_loop_intf_13.cur_state = AESL_inst_master.grp_convolution2_fu_344.ap_CS_fsm;
    assign seq_loop_intf_13.iter_start_state = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state5;
    assign seq_loop_intf_13.iter_end_state0 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state12;
    assign seq_loop_intf_13.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_13.one_state_loop = 1'b0;
    assign seq_loop_intf_13.one_state_block = 1'b0;
    assign seq_loop_intf_13.finish = finish;
    csv_file_dump seq_loop_csv_dumper_13;
    seq_loop_monitor #(42) seq_loop_monitor_13;
    seq_loop_intf#(42) seq_loop_intf_14(clock,reset);
    assign seq_loop_intf_14.pre_loop_state0 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state5;
    assign seq_loop_intf_14.pre_states_valid = 1'b1;
    assign seq_loop_intf_14.post_loop_state0 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state41;
    assign seq_loop_intf_14.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_14.post_loop_state1 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state21;
    assign seq_loop_intf_14.post_states_valid[1] = 1'b1;
    assign seq_loop_intf_14.post_loop_state2 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state29;
    assign seq_loop_intf_14.post_states_valid[2] = 1'b1;
    assign seq_loop_intf_14.quit_loop_state0 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state13;
    assign seq_loop_intf_14.quit_states_valid = 1'b1;
    assign seq_loop_intf_14.cur_state = AESL_inst_master.grp_convolution2_fu_344.ap_CS_fsm;
    assign seq_loop_intf_14.iter_start_state = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state13;
    assign seq_loop_intf_14.iter_end_state0 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state20;
    assign seq_loop_intf_14.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_14.one_state_loop = 1'b0;
    assign seq_loop_intf_14.one_state_block = 1'b0;
    assign seq_loop_intf_14.finish = finish;
    csv_file_dump seq_loop_csv_dumper_14;
    seq_loop_monitor #(42) seq_loop_monitor_14;
    seq_loop_intf#(42) seq_loop_intf_15(clock,reset);
    assign seq_loop_intf_15.pre_loop_state0 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state13;
    assign seq_loop_intf_15.pre_states_valid = 1'b1;
    assign seq_loop_intf_15.post_loop_state0 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state41;
    assign seq_loop_intf_15.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_15.post_loop_state1 = 42'h0;
    assign seq_loop_intf_15.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_15.post_loop_state2 = 42'h0;
    assign seq_loop_intf_15.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_15.quit_loop_state0 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state29;
    assign seq_loop_intf_15.quit_states_valid = 1'b1;
    assign seq_loop_intf_15.cur_state = AESL_inst_master.grp_convolution2_fu_344.ap_CS_fsm;
    assign seq_loop_intf_15.iter_start_state = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state29;
    assign seq_loop_intf_15.iter_end_state0 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state40;
    assign seq_loop_intf_15.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_15.one_state_loop = 1'b0;
    assign seq_loop_intf_15.one_state_block = 1'b0;
    assign seq_loop_intf_15.finish = finish;
    csv_file_dump seq_loop_csv_dumper_15;
    seq_loop_monitor #(42) seq_loop_monitor_15;
    seq_loop_intf#(42) seq_loop_intf_16(clock,reset);
    assign seq_loop_intf_16.pre_loop_state0 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state13;
    assign seq_loop_intf_16.pre_states_valid = 1'b1;
    assign seq_loop_intf_16.post_loop_state0 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state41;
    assign seq_loop_intf_16.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_16.post_loop_state1 = 42'h0;
    assign seq_loop_intf_16.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_16.post_loop_state2 = 42'h0;
    assign seq_loop_intf_16.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_16.quit_loop_state0 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state21;
    assign seq_loop_intf_16.quit_states_valid = 1'b1;
    assign seq_loop_intf_16.cur_state = AESL_inst_master.grp_convolution2_fu_344.ap_CS_fsm;
    assign seq_loop_intf_16.iter_start_state = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state21;
    assign seq_loop_intf_16.iter_end_state0 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state28;
    assign seq_loop_intf_16.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_16.one_state_loop = 1'b0;
    assign seq_loop_intf_16.one_state_block = 1'b0;
    assign seq_loop_intf_16.finish = finish;
    csv_file_dump seq_loop_csv_dumper_16;
    seq_loop_monitor #(42) seq_loop_monitor_16;
    seq_loop_intf#(42) seq_loop_intf_17(clock,reset);
    assign seq_loop_intf_17.pre_loop_state0 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state3;
    assign seq_loop_intf_17.pre_states_valid = 1'b1;
    assign seq_loop_intf_17.post_loop_state0 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state2;
    assign seq_loop_intf_17.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_17.post_loop_state1 = 42'h0;
    assign seq_loop_intf_17.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_17.post_loop_state2 = 42'h0;
    assign seq_loop_intf_17.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_17.quit_loop_state0 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state4;
    assign seq_loop_intf_17.quit_states_valid = 1'b1;
    assign seq_loop_intf_17.cur_state = AESL_inst_master.grp_convolution2_fu_344.ap_CS_fsm;
    assign seq_loop_intf_17.iter_start_state = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state4;
    assign seq_loop_intf_17.iter_end_state0 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state42;
    assign seq_loop_intf_17.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_17.one_state_loop = 1'b0;
    assign seq_loop_intf_17.one_state_block = 1'b0;
    assign seq_loop_intf_17.finish = finish;
    csv_file_dump seq_loop_csv_dumper_17;
    seq_loop_monitor #(42) seq_loop_monitor_17;
    seq_loop_intf#(42) seq_loop_intf_18(clock,reset);
    assign seq_loop_intf_18.pre_loop_state0 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state1;
    assign seq_loop_intf_18.pre_states_valid = 1'b1;
    assign seq_loop_intf_18.post_loop_state0 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state1;
    assign seq_loop_intf_18.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_18.post_loop_state1 = 42'h0;
    assign seq_loop_intf_18.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_18.post_loop_state2 = 42'h0;
    assign seq_loop_intf_18.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_18.quit_loop_state0 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state2;
    assign seq_loop_intf_18.quit_states_valid = 1'b1;
    assign seq_loop_intf_18.cur_state = AESL_inst_master.grp_convolution2_fu_344.ap_CS_fsm;
    assign seq_loop_intf_18.iter_start_state = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state2;
    assign seq_loop_intf_18.iter_end_state0 = AESL_inst_master.grp_convolution2_fu_344.ap_ST_fsm_state4;
    assign seq_loop_intf_18.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_18.one_state_loop = 1'b0;
    assign seq_loop_intf_18.one_state_block = 1'b0;
    assign seq_loop_intf_18.finish = finish;
    csv_file_dump seq_loop_csv_dumper_18;
    seq_loop_monitor #(42) seq_loop_monitor_18;
    seq_loop_intf#(9) seq_loop_intf_19(clock,reset);
    assign seq_loop_intf_19.pre_loop_state0 = AESL_inst_master.grp_maxPool_fu_354.ap_ST_fsm_state5;
    assign seq_loop_intf_19.pre_states_valid = 1'b1;
    assign seq_loop_intf_19.post_loop_state0 = AESL_inst_master.grp_maxPool_fu_354.ap_ST_fsm_state3;
    assign seq_loop_intf_19.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_19.post_loop_state1 = 9'h0;
    assign seq_loop_intf_19.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_19.post_loop_state2 = 9'h0;
    assign seq_loop_intf_19.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_19.quit_loop_state0 = AESL_inst_master.grp_maxPool_fu_354.ap_ST_fsm_state6;
    assign seq_loop_intf_19.quit_states_valid = 1'b1;
    assign seq_loop_intf_19.cur_state = AESL_inst_master.grp_maxPool_fu_354.ap_CS_fsm;
    assign seq_loop_intf_19.iter_start_state = AESL_inst_master.grp_maxPool_fu_354.ap_ST_fsm_state6;
    assign seq_loop_intf_19.iter_end_state0 = AESL_inst_master.grp_maxPool_fu_354.ap_ST_fsm_state9;
    assign seq_loop_intf_19.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_19.one_state_loop = 1'b0;
    assign seq_loop_intf_19.one_state_block = 1'b0;
    assign seq_loop_intf_19.finish = finish;
    csv_file_dump seq_loop_csv_dumper_19;
    seq_loop_monitor #(9) seq_loop_monitor_19;
    seq_loop_intf#(9) seq_loop_intf_20(clock,reset);
    assign seq_loop_intf_20.pre_loop_state0 = AESL_inst_master.grp_maxPool_fu_354.ap_ST_fsm_state2;
    assign seq_loop_intf_20.pre_states_valid = 1'b1;
    assign seq_loop_intf_20.post_loop_state0 = AESL_inst_master.grp_maxPool_fu_354.ap_ST_fsm_state2;
    assign seq_loop_intf_20.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_20.post_loop_state1 = 9'h0;
    assign seq_loop_intf_20.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_20.post_loop_state2 = 9'h0;
    assign seq_loop_intf_20.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_20.quit_loop_state0 = AESL_inst_master.grp_maxPool_fu_354.ap_ST_fsm_state3;
    assign seq_loop_intf_20.quit_states_valid = 1'b1;
    assign seq_loop_intf_20.cur_state = AESL_inst_master.grp_maxPool_fu_354.ap_CS_fsm;
    assign seq_loop_intf_20.iter_start_state = AESL_inst_master.grp_maxPool_fu_354.ap_ST_fsm_state3;
    assign seq_loop_intf_20.iter_end_state0 = AESL_inst_master.grp_maxPool_fu_354.ap_ST_fsm_state6;
    assign seq_loop_intf_20.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_20.one_state_loop = 1'b0;
    assign seq_loop_intf_20.one_state_block = 1'b0;
    assign seq_loop_intf_20.finish = finish;
    csv_file_dump seq_loop_csv_dumper_20;
    seq_loop_monitor #(9) seq_loop_monitor_20;
    seq_loop_intf#(9) seq_loop_intf_21(clock,reset);
    assign seq_loop_intf_21.pre_loop_state0 = AESL_inst_master.grp_maxPool_fu_354.ap_ST_fsm_state1;
    assign seq_loop_intf_21.pre_states_valid = 1'b1;
    assign seq_loop_intf_21.post_loop_state0 = AESL_inst_master.grp_maxPool_fu_354.ap_ST_fsm_state1;
    assign seq_loop_intf_21.post_states_valid[0] = 1'b1;
    assign seq_loop_intf_21.post_loop_state1 = 9'h0;
    assign seq_loop_intf_21.post_states_valid[1] = 1'b0;
    assign seq_loop_intf_21.post_loop_state2 = 9'h0;
    assign seq_loop_intf_21.post_states_valid[2] = 1'b0;
    assign seq_loop_intf_21.quit_loop_state0 = AESL_inst_master.grp_maxPool_fu_354.ap_ST_fsm_state2;
    assign seq_loop_intf_21.quit_states_valid = 1'b1;
    assign seq_loop_intf_21.cur_state = AESL_inst_master.grp_maxPool_fu_354.ap_CS_fsm;
    assign seq_loop_intf_21.iter_start_state = AESL_inst_master.grp_maxPool_fu_354.ap_ST_fsm_state2;
    assign seq_loop_intf_21.iter_end_state0 = AESL_inst_master.grp_maxPool_fu_354.ap_ST_fsm_state3;
    assign seq_loop_intf_21.iter_end_states_valid = 1'b1;
    assign seq_loop_intf_21.one_state_loop = 1'b0;
    assign seq_loop_intf_21.one_state_block = 1'b0;
    assign seq_loop_intf_21.finish = finish;
    csv_file_dump seq_loop_csv_dumper_21;
    seq_loop_monitor #(9) seq_loop_monitor_21;
    upc_loop_intf#(1) upc_loop_intf_1(clock,reset);
    assign upc_loop_intf_1.cur_state = AESL_inst_master.grp_master_Pipeline_VITIS_LOOP_143_2_fu_360.ap_CS_fsm;
    assign upc_loop_intf_1.iter_start_state = AESL_inst_master.grp_master_Pipeline_VITIS_LOOP_143_2_fu_360.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_end_state = AESL_inst_master.grp_master_Pipeline_VITIS_LOOP_143_2_fu_360.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.quit_state = AESL_inst_master.grp_master_Pipeline_VITIS_LOOP_143_2_fu_360.ap_ST_fsm_pp0_stage0;
    assign upc_loop_intf_1.iter_start_block = AESL_inst_master.grp_master_Pipeline_VITIS_LOOP_143_2_fu_360.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_end_block = AESL_inst_master.grp_master_Pipeline_VITIS_LOOP_143_2_fu_360.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.quit_block = AESL_inst_master.grp_master_Pipeline_VITIS_LOOP_143_2_fu_360.ap_block_pp0_stage0_subdone;
    assign upc_loop_intf_1.iter_start_enable = AESL_inst_master.grp_master_Pipeline_VITIS_LOOP_143_2_fu_360.ap_enable_reg_pp0_iter0;
    assign upc_loop_intf_1.iter_end_enable = AESL_inst_master.grp_master_Pipeline_VITIS_LOOP_143_2_fu_360.ap_enable_reg_pp0_iter31;
    assign upc_loop_intf_1.quit_enable = AESL_inst_master.grp_master_Pipeline_VITIS_LOOP_143_2_fu_360.ap_enable_reg_pp0_iter31;
    assign upc_loop_intf_1.loop_start = AESL_inst_master.grp_master_Pipeline_VITIS_LOOP_143_2_fu_360.ap_start;
    assign upc_loop_intf_1.loop_ready = AESL_inst_master.grp_master_Pipeline_VITIS_LOOP_143_2_fu_360.ap_ready;
    assign upc_loop_intf_1.loop_done = AESL_inst_master.grp_master_Pipeline_VITIS_LOOP_143_2_fu_360.ap_done_int;
    assign upc_loop_intf_1.loop_continue = 1'b1;
    assign upc_loop_intf_1.quit_at_end = 1'b1;
    assign upc_loop_intf_1.finish = finish;
    csv_file_dump upc_loop_csv_dumper_1;
    upc_loop_monitor #(1) upc_loop_monitor_1;

    sample_manager sample_manager_inst;

initial begin
    sample_manager_inst = new;



    mstatus_csv_dumper_1 = new("./module_status1.csv");
    module_monitor_1 = new(module_intf_1,mstatus_csv_dumper_1);
    mstatus_csv_dumper_2 = new("./module_status2.csv");
    module_monitor_2 = new(module_intf_2,mstatus_csv_dumper_2);
    mstatus_csv_dumper_3 = new("./module_status3.csv");
    module_monitor_3 = new(module_intf_3,mstatus_csv_dumper_3);
    mstatus_csv_dumper_4 = new("./module_status4.csv");
    module_monitor_4 = new(module_intf_4,mstatus_csv_dumper_4);
    mstatus_csv_dumper_5 = new("./module_status5.csv");
    module_monitor_5 = new(module_intf_5,mstatus_csv_dumper_5);
    mstatus_csv_dumper_6 = new("./module_status6.csv");
    module_monitor_6 = new(module_intf_6,mstatus_csv_dumper_6);



    seq_loop_csv_dumper_1 = new("./seq_loop_status1.csv");
    seq_loop_monitor_1 = new(seq_loop_intf_1,seq_loop_csv_dumper_1);
    seq_loop_csv_dumper_2 = new("./seq_loop_status2.csv");
    seq_loop_monitor_2 = new(seq_loop_intf_2,seq_loop_csv_dumper_2);
    seq_loop_csv_dumper_3 = new("./seq_loop_status3.csv");
    seq_loop_monitor_3 = new(seq_loop_intf_3,seq_loop_csv_dumper_3);
    seq_loop_csv_dumper_4 = new("./seq_loop_status4.csv");
    seq_loop_monitor_4 = new(seq_loop_intf_4,seq_loop_csv_dumper_4);
    seq_loop_csv_dumper_5 = new("./seq_loop_status5.csv");
    seq_loop_monitor_5 = new(seq_loop_intf_5,seq_loop_csv_dumper_5);
    seq_loop_csv_dumper_6 = new("./seq_loop_status6.csv");
    seq_loop_monitor_6 = new(seq_loop_intf_6,seq_loop_csv_dumper_6);
    seq_loop_csv_dumper_7 = new("./seq_loop_status7.csv");
    seq_loop_monitor_7 = new(seq_loop_intf_7,seq_loop_csv_dumper_7);
    seq_loop_csv_dumper_8 = new("./seq_loop_status8.csv");
    seq_loop_monitor_8 = new(seq_loop_intf_8,seq_loop_csv_dumper_8);
    seq_loop_csv_dumper_9 = new("./seq_loop_status9.csv");
    seq_loop_monitor_9 = new(seq_loop_intf_9,seq_loop_csv_dumper_9);
    seq_loop_csv_dumper_10 = new("./seq_loop_status10.csv");
    seq_loop_monitor_10 = new(seq_loop_intf_10,seq_loop_csv_dumper_10);
    seq_loop_csv_dumper_11 = new("./seq_loop_status11.csv");
    seq_loop_monitor_11 = new(seq_loop_intf_11,seq_loop_csv_dumper_11);
    seq_loop_csv_dumper_12 = new("./seq_loop_status12.csv");
    seq_loop_monitor_12 = new(seq_loop_intf_12,seq_loop_csv_dumper_12);
    seq_loop_csv_dumper_13 = new("./seq_loop_status13.csv");
    seq_loop_monitor_13 = new(seq_loop_intf_13,seq_loop_csv_dumper_13);
    seq_loop_csv_dumper_14 = new("./seq_loop_status14.csv");
    seq_loop_monitor_14 = new(seq_loop_intf_14,seq_loop_csv_dumper_14);
    seq_loop_csv_dumper_15 = new("./seq_loop_status15.csv");
    seq_loop_monitor_15 = new(seq_loop_intf_15,seq_loop_csv_dumper_15);
    seq_loop_csv_dumper_16 = new("./seq_loop_status16.csv");
    seq_loop_monitor_16 = new(seq_loop_intf_16,seq_loop_csv_dumper_16);
    seq_loop_csv_dumper_17 = new("./seq_loop_status17.csv");
    seq_loop_monitor_17 = new(seq_loop_intf_17,seq_loop_csv_dumper_17);
    seq_loop_csv_dumper_18 = new("./seq_loop_status18.csv");
    seq_loop_monitor_18 = new(seq_loop_intf_18,seq_loop_csv_dumper_18);
    seq_loop_csv_dumper_19 = new("./seq_loop_status19.csv");
    seq_loop_monitor_19 = new(seq_loop_intf_19,seq_loop_csv_dumper_19);
    seq_loop_csv_dumper_20 = new("./seq_loop_status20.csv");
    seq_loop_monitor_20 = new(seq_loop_intf_20,seq_loop_csv_dumper_20);
    seq_loop_csv_dumper_21 = new("./seq_loop_status21.csv");
    seq_loop_monitor_21 = new(seq_loop_intf_21,seq_loop_csv_dumper_21);

    upc_loop_csv_dumper_1 = new("./upc_loop_status1.csv");
    upc_loop_monitor_1 = new(upc_loop_intf_1,upc_loop_csv_dumper_1);

    sample_manager_inst.add_one_monitor(module_monitor_1);
    sample_manager_inst.add_one_monitor(module_monitor_2);
    sample_manager_inst.add_one_monitor(module_monitor_3);
    sample_manager_inst.add_one_monitor(module_monitor_4);
    sample_manager_inst.add_one_monitor(module_monitor_5);
    sample_manager_inst.add_one_monitor(module_monitor_6);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_1);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_2);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_3);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_4);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_5);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_6);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_7);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_8);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_9);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_10);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_11);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_12);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_13);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_14);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_15);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_16);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_17);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_18);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_19);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_20);
    sample_manager_inst.add_one_monitor(seq_loop_monitor_21);
    sample_manager_inst.add_one_monitor(upc_loop_monitor_1);
    
    fork
        sample_manager_inst.start_monitor();
        last_transaction_done;
    join
    disable fork;

    sample_manager_inst.start_dump();
end

    task last_transaction_done();
        wait(reset == 0);
        while(1) begin
            if (finish == 1'b1)
                break;
            else
                @(posedge clock);
        end
    endtask


endmodule
